always_ff @